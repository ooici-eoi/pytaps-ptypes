test_data/roms.nc.cdl