test_data/coads.nc.cdl