test_data/ncom.nc.cdl