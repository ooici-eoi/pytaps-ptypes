test_data/usgs.nc.cdl