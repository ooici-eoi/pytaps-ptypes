book    mark    8   8   4�           �R��0��A       T�       Users        cmueller     Development      OOI      Dev 	     datamodel        pytaps-ptypes   	     test_data   
     hfr.nc.cdl  $           $   8   D   P   d   |   �        �:          S�          �	          ��+          ��+          �Ή          q��          ���          '��     $     �   �   �           0  @  P                                         �       Macintosh HD      �?Tt         A���   $     6D95C714-29C8-30BC-A452-DE34B50798C2     �     �?                 /                 �    icns  �is32  ���� ��  ��� �� ��ߥ� �� ����� �� ������� �� ������ �� ������� �� ����� �� ���� �� ���� �� ���� �� ���� �� ���� ��  ��  ��  ��  ��� ����� ��  ��� �� ��ߥ� �� ����� �� ������� �� ������ �� ������� �� ����� �� ���� �� ���� �� ���� �� ���� �� ���� ��  ��  ��  ��  ��� ����� ��  ��� �� ��ߥ� �� ����� �� ������� �� ������ �� ������� �� ����� �� ���� �� ���� �� ���� �� ���� �� ���� ��  ��  ��  ��  ��� ��s8mk    +8888888        8�������8       9��������9      9���������9     :����������:    ;����������;    =����������=    >����������>    ?����������?    @����������@    A����������A    C����������C    D����������D    E����������E    E����������E    6OXdknnkdXO6  il32  ܁�� ��  �������X� �� �����ʴ�S� �� ����Ь��Q� �� ����ֵ���N� �� ����������M� �� ����˥����L� �� ����ӧ�����J  �� ��
�ڷ}a_k��D �� ��	�ӻ������ �� ������ĳ�� �� �������ʿ� �� ��������� �� �������� �� ������� �� ������� �� ����� �� ������ �� ����� �� ���� �� ���� �� ���� �� ���� �� ���� �� ���� �� ���� �� ���� �� ���� �� ���� ��  ��  ��� ��� ����� ��  �������X� �� �����ʴ�S� �� ����Ь��Q� �� ����ֵ���N� �� ����������M� �� ����˥����L� �� ����ӧ�����J  �� ��
�ڷ}a_k��D �� ��	�ӻ������ �� ������ĳ�� �� �������ʿ� �� ��������� �� �������� �� ������� �� ������� �� ����� �� ������ �� ����� �� ���� �� ���� �� ���� �� ���� �� ���� �� ���� �� ���� �� ���� �� ���� �� ���� ��  ��  ��� ��� ����� ��  �������X� �� �����ʴ�S� �� ����Ь��Q� �� ����ֵ���N� �� ����������M� �� ����˥����L� �� ����ӧ�����J  �� ��
�ڷ}a_k��D �� ��	�ӻ������ �� ������ĳ�� �� �������ʿ� �� ��������� �� �������� �� ������� �� ������� �� ����� �� ������ �� ����� �� ���� �� ���� �� ���� �� ���� �� ���� �� ���� �� ���� �� ���� �� ���� �� ���� ��  ��  ��� ��� ��l8mk      -MMMMMMMMMMMMM?                M��������������m                O���������������r               T����������������r              V�����������������s             V������������������s            V�������������������s           V��������������������s          V���������������������m         V����������������������@        V����������������������P        V����������������������S        V����������������������U        V����������������������V        V����������������������V        V����������������������V        V����������������������V        V����������������������V        V����������������������V        V����������������������V        V����������������������V        V����������������������V        V����������������������V        V����������������������V        V����������������������V        V����������������������V        V����������������������V        V����������������������V        V����������������������V        V����������������������V        8dmmmmmmmmmmmmmmmmmmmmd8        
!!!!!!!!!!!!!!!!!!!!
    it32      ��� ��� ��� ��������Ӥ0� ��� ��� ���������������1� ��� ��� �����	���������h� ��� ��� �����������������o� ��� ��� ��������������ƿ�d� ��� ��� ����������������Ľ��b� ��� ��� ���������������Ľ���a� ��� ��� ���������������Ľ����`� ��� ��� ���������������ƽ�����`� ��� ��� ���������������������`� ��� ��� ���������������ĺ������`� ��� ��� ��������������Ǽ�������`� ��� ��� ����������������������_� ��� ��� ��������������ĸ��������_� ��� ��� �������������ź���������_� ��� ��� ������������ƻ����������`� ��� ��� ������������ɾ�����������`� ��� ��� �����������˿������������b� ��� ��� ��������������������������a� ��� ��� �����������µ�������������c� ��� ��� �����������¶��������������c� ��� ��� �����������÷����
����������d� ��� ��� �����������Ź����
����������d� ��� ��� �����������ƻ����
����������f� ��� ��� �����������Ǽ���
����������h� ��� ��� �����������ɿ�������������������h� ��� ��� �����������������}wtrpnlr��������h�  �� ��� �� ����������¸����}{{yxwtsqoko����d� ��� ������������ż�������~|�zyywqw��V� ��� ����������������������������|u��7� ��� �������������û������������������{�� ��� ��"������������������������������������ ��� ������������������������������������G� ��� ���������������ÿ�������������������� ��� ��#������������������������������������� ��� �����������������́� ʁ�	����������� ��� �������������������т������������́ ��� ����������������ډ�������Ձ ��� �������������������߃�������ہ ��� ������������������������� ��� ������������	���������� ��� ���������� � ��� �������� � ��� ������ � ��� ����� ��� ���� ��� ���� ��� �� ��� �� ��� �� ��� �� ��� �� ��� �� ��� �� ��� �� ��� �� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��������� ��� ��� ��������Ӥ0� ��� ��� ���������������1� ��� ��� �����	���������h� ��� ��� �����������������o� ��� ��� ��������������ƿ�d� ��� ��� ����������������Ľ��b� ��� ��� ���������������Ľ���a� ��� ��� ���������������Ľ����`� ��� ��� ���������������ƽ�����`� ��� ��� ���������������������`� ��� ��� ���������������ĺ������`� ��� ��� ��������������Ǽ�������`� ��� ��� ����������������������_� ��� ��� ��������������ĸ��������_� ��� ��� �������������ź���������_� ��� ��� ������������ƻ����������`� ��� ��� ������������ɾ�����������`� ��� ��� �����������˿������������b� ��� ��� ��������������������������a� ��� ��� �����������µ�������������c� ��� ��� �����������¶��������������c� ��� ��� �����������÷����
����������d� ��� ��� �����������Ź����
����������d� ��� ��� �����������ƻ����
����������f� ��� ��� �����������Ǽ���
����������h� ��� ��� �����������ɿ�������������������h� ��� ��� �����������������}wtrpnlr��������h�  �� ��� �� ����������¸����}{{yxwtsqoko����d� ��� ������������ż�������~|�zyywqw��V� ��� ����������������������������|u��7� ��� �������������û������������������{�� ��� ��"������������������������������������ ��� ������������������������������������G� ��� ���������������ÿ�������������������� ��� ��#������������������������������������� ��� �����������������́� ʁ�	����������� ��� �������������������т������������́ ��� ����������������ډ�������Ձ ��� �������������������߃�������ہ ��� ������������������������� ��� ������������	���������� ��� ���������� � ��� �������� � ��� ������ � ��� ����� ��� ���� ��� ���� ��� �� ��� �� ��� �� ��� �� ��� �� ��� �� ��� �� ��� �� ��� �� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��������� ��� ��� ��������Ӥ0� ��� ��� ���������������1� ��� ��� �����	���������h� ��� ��� �����������������o� ��� ��� ��������������ƿ�d� ��� ��� ����������������Ľ��b� ��� ��� ���������������Ľ���a� ��� ��� ���������������Ľ����`� ��� ��� ���������������ƽ�����`� ��� ��� ���������������������`� ��� ��� ���������������ĺ������`� ��� ��� ��������������Ǽ�������`� ��� ��� ����������������������_� ��� ��� ��������������ĸ��������_� ��� ��� �������������ź���������_� ��� ��� ������������ƻ����������`� ��� ��� ������������ɾ�����������`� ��� ��� �����������˿������������b� ��� ��� ��������������������������a� ��� ��� �����������µ�������������c� ��� ��� �����������¶��������������c� ��� ��� �����������÷����
����������d� ��� ��� �����������Ź����
����������d� ��� ��� �����������ƻ����
����������f� ��� ��� �����������Ǽ���
����������h� ��� ��� �����������ɿ�������������������h� ��� ��� �����������������}wtrpnlr��������h�  �� ��� �� ����������¸����}{{yxwtsqoko����d� ��� ������������ż�������~|�zyywqw��V� ��� ����������������������������|u��7� ��� �������������û������������������{�� ��� ��"������������������������������������ ��� ������������������������������������G� ��� ���������������ÿ�������������������� ��� ��#������������������������������������� ��� �����������������́� ʁ�	����������� ��� �������������������т������������́ ��� ����������������ډ�������Ձ ��� �������������������߃�������ہ ��� ������������������������� ��� ������������	���������� ��� ���������� � ��� �������� � ��� ������ � ��� ����� ��� ���� ��� ���� ��� �� ��� �� ��� �� ��� �� ��� �� ��� �� ��� �� ��� �� ��� �� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ������t8mk  @                                                                                 +012222222222222222222222222222222222222222222222221/+#
                                                              	�������������������������������������������������������u;                                                             *�����������������������������������������������������������8                                                            3������������������������������������������������������������W                                                           <�������������������������������������������������������������^                                                           C��������������������������������������������������������������Z                                                         "E���������������������������������������������������������������V                                                        $G����������������������������������������������������������������S                                                       $G�����������������������������������������������������������������S                                                      $G������������������������������������������������������������������R                                                     $G�������������������������������������������������������������������R                                                    $G��������������������������������������������������������������������R                                                   $G���������������������������������������������������������������������Q                                                  $G����������������������������������������������������������������������R                                                 $G�����������������������������������������������������������������������R                                                $G������������������������������������������������������������������������R                                               $F�������������������������������������������������������������������������Q                                              $F��������������������������������������������������������������������������Q                                             $F���������������������������������������������������������������������������P                                            $E����������������������������������������������������������������������������Q                                           $E�����������������������������������������������������������������������������P                                          $E������������������������������������������������������������������������������P                                         $E�������������������������������������������������������������������������������P                                        $E��������������������������������������������������������������������������������P                                       $E���������������������������������������������������������������������������������O                                      $E����������������������������������������������������������������������������������N                                     $E�����������������������������������������������������������������������������������N                                    $E������������������������������������������������������������������������������������L                                   $E�������������������������������������������������������������������������������������J                                  $D��������������������������������������������������������������������������������������E                                 $D���������������������������������������������������������������������������������������:                                $D����������������������������������������������������������������������������������������)                               $C�����������������������������������������������������������������������������������������                               $C�����������������������������������������������������������������������������������������?                              $C������������������������������������������������������������������������������������������                               $B������������������������������������������������������������������������������������������,                              $B������������������������������������������������������������������������������������������6	                              $B������������������������������������������������������������������������������������������<                              $B������������������������������������������������������������������������������������������A                              $B������������������������������������������������������������������������������������������D                               $B������������������������������������������������������������������������������������������E"                              $B������������������������������������������������������������������������������������������E"                              $A������������������������������������������������������������������������������������������E#                              $A������������������������������������������������������������������������������������������E#                              $A������������������������������������������������������������������������������������������E#                              $A������������������������������������������������������������������������������������������E#                              $@������������������������������������������������������������������������������������������E#                              $@������������������������������������������������������������������������������������������E$                              $@������������������������������������������������������������������������������������������E$                              $@������������������������������������������������������������������������������������������E$                              $@������������������������������������������������������������������������������������������E$                              $@������������������������������������������������������������������������������������������E$                              $@������������������������������������������������������������������������������������������E$                              $@������������������������������������������������������������������������������������������E$                              $@������������������������������������������������������������������������������������������E$                              $@������������������������������������������������������������������������������������������E$                              $@������������������������������������������������������������������������������������������E$                              $?������������������������������������������������������������������������������������������E$                              $?������������������������������������������������������������������������������������������E$                              $?������������������������������������������������������������������������������������������E$                              $?������������������������������������������������������������������������������������������D$                              $?������������������������������������������������������������������������������������������D$                              $?������������������������������������������������������������������������������������������D$                              $?������������������������������������������������������������������������������������������D$                              $?������������������������������������������������������������������������������������������C$                              $?������������������������������������������������������������������������������������������C$                              $?������������������������������������������������������������������������������������������C$                              $?������������������������������������������������������������������������������������������C$                              $?������������������������������������������������������������������������������������������C$                              $?������������������������������������������������������������������������������������������C$                              $?������������������������������������������������������������������������������������������B$                              $?������������������������������������������������������������������������������������������B$                              $?������������������������������������������������������������������������������������������B$                              $?������������������������������������������������������������������������������������������B$                              $?������������������������������������������������������������������������������������������B$                              $?������������������������������������������������������������������������������������������B$                              $?������������������������������������������������������������������������������������������B$                              $>������������������������������������������������������������������������������������������B$                              $>������������������������������������������������������������������������������������������B$                              $>������������������������������������������������������������������������������������������B$                              $>������������������������������������������������������������������������������������������A$                              $>������������������������������������������������������������������������������������������A$                              $>������������������������������������������������������������������������������������������A$                              $>������������������������������������������������������������������������������������������A$                              $>������������������������������������������������������������������������������������������A$                              $>������������������������������������������������������������������������������������������A$                              $>������������������������������������������������������������������������������������������A$                              $>������������������������������������������������������������������������������������������@$                              $>������������������������������������������������������������������������������������������@$                              $=������������������������������������������������������������������������������������������@$                              $=������������������������������������������������������������������������������������������@$                              $=������������������������������������������������������������������������������������������@$                              $=������������������������������������������������������������������������������������������@$                              $=������������������������������������������������������������������������������������������@$                              $=������������������������������������������������������������������������������������������?$                              $=������������������������������������������������������������������������������������������?$                              $=������������������������������������������������������������������������������������������?$                              $=������������������������������������������������������������������������������������������?$                              $=������������������������������������������������������������������������������������������?$                              $=������������������������������������������������������������������������������������������?$                              $=������������������������������������������������������������������������������������������?$                              $=������������������������������������������������������������������������������������������?$                              $=������������������������������������������������������������������������������������������?$                              $=������������������������������������������������������������������������������������������?$                              $=������������������������������������������������������������������������������������������?$                              $<������������������������������������������������������������������������������������������?$                              $<������������������������������������������������������������������������������������������?$                              $<������������������������������������������������������������������������������������������?$                              $<������������������������������������������������������������������������������������������?$                              $<������������������������������������������������������������������������������������������?$                              $<������������������������������������������������������������������������������������������>$                              $<������������������������������������������������������������������������������������������>$                              $<������������������������������������������������������������������������������������������>$                              $<������������������������������������������������������������������������������������������>$                              $<������������������������������������������������������������������������������������������>$                              $<������������������������������������������������������������������������������������������>$                              $<������������������������������������������������������������������������������������������>$                              ";������������������������������������������������������������������������������������������<"                               6������������������������������������������������������������������������������������������7                               .EWenssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssofXF/                              $6EOWZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZWOE6$                              $.5:<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<:5.$                              	 "$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$" 	                                                                                                                                                                                                                                                                                                                                             ic08  k   jP  
�
   ftypjp2     jp2    Ojp2h   ihdr           colr        "cdef                      jp2c�O�Q 2                               �R     �\  PXX`XX`XX`XXXPPX�d  Kakadu-v5.2.1�� 
    ~ ����o�D���Ht�����0��_ꏓ�q6e!V	�1q�4�� }3:f!�@T$������f� ����� _�Wt8�yL��X)c,/ʲ��V6Bh|r��f�1,Ŀ��B��6�v�o���~�����P���]�D? 5L,ZS{2L���Kj ��ia���0�(�x�6�V���n�Jٟ�+H��⏃��O�_��1�����7�'�؜xK7[�|:X�'+3�0�56��"�̂���F?
A~�aj��p�倀��I��~c@�����?��T��k�"~�&
�9�`���٠����<����Ip��~�]���gK�Ј��;�/��+��Ia�̂!�@�;c6��=C����~h ��c���	۫~�$�����6G���;���	�B�b2�����U*�2
��S)�m�
z�F4�Wݻ?��(�Ӏ����H��X�l(�����eo���*K@����(�6��J�_���eat:-u�"6
� hC��

��g�����&L�@%� ��D��=�!܎� �<^5Q$8��ܠ����F��2��u�E��w��ϒ��S��>ᎌ�5"���R��=_�]���'!.��b?e�7T����vK^��������?���θ�M�]����*F�*�3R�N�J�%
A�n5~�_���]��7�U#��_G�p#�q�ӌ�D�J�N𓚉,�5�"c�������Of���"�"D:�����أU߸�8�����	������z��A�꾪��5�.?<��w�ƋN�ds�C���Q7����̻<b3G��۟���؆��3�.bq�R-_�@���S��UD'R�a�b�k����^��/=%�SÑ��y�D�qyo��;����#�'��|"���Ny����4��1��H� H����)�|�R\���[Р��K ����4b�Z��|4LqЀ�M޾������ӟJ�i��$�y�X�ڲZ5$��V�LN�$�P�q7��P�7'����lW�4�O���i�%�#��Nh��K��B�~�A����   )=L_D��kB<d��ȇ�ҥ)J'�J�2�-�'�������(�j���y�pl�q�RE��*� ����w��]E/����ےI$�fr��R��b,����AB��l�% ���I$�I$�t��K�EGMC��[E�W�2���b\�V��f�`���gg���Ҥ��7Zƨ����^��jQw`�o�e�����g�����z��������?�Ņ��6�G�t��	`g����@�����u�E	�(�v�M&��@1)������Q @SC]�-lHMV���@�p��l k�߁؁��8<-t���w����@C�h��p¶�q������w� /vZ��{�&A�-��[u����w�w�D	-W  ,�� �oh�p��Ǻ��SvF:#.X���w��WW��)!&�`z3�����S���\��)�
3�5���r��$����R�'a,��m�K�F`{��:R�2�E��n� �g��Tԣ<�^�jZ[��a Cq"ㅐ��a@  ĝYjGw��\�"  ����\��P�6��xT�πw`�o�Q
n�R�-��4�?8����ҽ>�}���p��ҁԖ����j|����2���s��x�.�5I�� �}��u|Ǩ���N,I�ǁ~9� J��즦A�pj��y���)��t2�ypĭr�do`K�o��F� ��`�-[����L%�$�4�[�Jˬ�sX���ixެ7����3,4ٮ���$��H��/)yKɳ Z�|�7��+���0�ݲ��AF�(8J�Iz�
��0B׎�yy��f�h��Z�0�raڰ��{>����oG�������J�6<���I�|�N1�ӈ�����P��D�so��c�!MK�wsӗ߇?�4��cjP��J�!��L	NWVI�a������"M<�fe+v��#B������G�֏ώ�ދ���7�{k��G�8��e)����:�7��6k�7�T��k��E���mQn�퐤�%�!�0p�e��]��L�-IC�u�E7�Y���D�b�b�)N��)�f������lD��E
�Ɍ:b3O�H��Xd��O/ϊ4�櫁`�u�9
~����k��m����[�r�oR֘84ݓ
_�E�$�k>)j��
<��S�N��x)�p�|�q�A��6���"M2:�Rv�p�B[
�f�W����T�]�%��sc��6�,���m�q�P����=u��-А#�A�s@$-��	�[��@[���6}]�^u�[\��f8�!�)�������Ԏ=m�/U�?
��BȈI    ��Lʠch
%(�N���:��)o�y֩��H�'�t4_��|�LH	�Z���(���>�$ZR7%�h$ !@h6�I$�I$�I$�I$�ڻE'��TL(0� t�ҩw��W��Wڶ�j�]��eM�~bb�	���\�k�"��މ҃�O��1d�M�����m�m�ິ�c�yA�$�I$�I$�I$�I>٧U�u�� �����B�B(��,#�O����Qy�փ�{��q#��.�f�l�Ky��q��W����o��xy�!_ӑj<��@cv��v2��9��<Uͽ �\�bn`U�/b�ړ��b�IED�u6�����5p���OgL*����&��&��4�ϻ���]��LNJቔc���'�4z1g�ۮ�C>��x��dׁ����4�+����nq�]�����S��zs���k?�e:�;��o��(Q<Ӷӏ�oQzZ<�O��	"�V���JT�6SK7��c/DE����#�#�[?��^Z��c�o�F#����ؖ�:\e��V�|�7��|��e.��"]E-�GA�j��f��??+ �(�Y�+�_7��|�7�z��t�F�T�d�FS�j�1,�7����?O���=��Ǎ5@�j��G��"%0\�S#T���������"�SLc����W��[�pe��_�W�J���L�!����Y���%��Gx��E��`Wأ��Ո�w��Au�o�OP0v�B�VP�E@C�`	,�q�7zA"�.�g�)���HNGU��o����y�f��=�u��F* �KR�/�l�Y%�e4�V�Cda�� h�6P�!p� 2���h�@Dd��]Q���#�vt�}��P  ���	D�\6��?,$%��A}�����_
Z�Qf�^*-�Q���N�!$�2�_�'(���D�K��f n�����.C��=Q:��Ad���s|�΄w���Q"
��W�!?���ڝ��3���<�����_h]���^R�D� `0�%�[e�#1EX��~�_7��|�7��|�7�v��N
(��$��_۴��u��{�V�G~i����x��kVr���癭?Ԙ��?+.l���]|�lU��b����I<������D�S�����
M�_�w'����B{�l�˟���s����:�r`��p��!�4�����M��j0G.��	}�oo��0�0��;
�{�3XYA꤉Z��ǔ�)�}���/IB�	�p�)�.�;Aku�~[���f}��Dܿ*�Ky�C0��h*���=M��ٛ}{�Hj� �F�>�x�OFf��_P��U����z�#
����n�n�9���)�cg��� D�
M�dX��F���&S��g�����*��=d�)z Xyl��k5�V�=l���p��}RwM��I�a�շ�u5:j�i��� �/K�+!��Ns�$,��IMg�b�VIV���?���	�U"P L6�gi�oK�l�3 � *>�۾U���l����r��HK2���/m����o:ݔK<���s^��b�ҟw�R\����#����W+o���Iڙ�!�=�K�������7�A .P�{�Fƀj8��X�9�� xI�����&r��Db�Y�J�︧g�(��l�]�*�^_�����H6��Q���p('�Hf�xD�b�����o����o�2,m���|�7��|�7��|�l� �q ��[u�|��'c�*�A�V�j��ET�:H�I�����O"+���@��b^��))b�P��$Q��X¶����o��?=P��[�#jtd/��c��V�|�d`�Z��}���l��8#�      6_�        �}P       {p��R�z������p)�:�^��'hл�&�c��z8No����!=�m���VV��ǫ�[�12��Ğ8 �6��P��W¿�Y�$�fш��R�� 0|�Ρv!:���yW��w�����  �U��?��   �STWt]|_���-è�g�VX���������1���H    Jڶ�An�tS�
���T�������BΝ�lWW\�     Y�zk?b��U�~a!�Jҁ��M�RuK���_��T �ٸ|[m��q�h�i:�A    o�i^̻gN����Lǆ�H##>���k�_���{k`��ډ���U��0��Y�Y����3�Z�D�((�Mogѻh+O���|�y-S��Rtc����''�-t"@��@��a�zdLD=<�����}�f۸8������f G�cP�;W�aU^�>�ZUF/���1W[�$ɚŨ4e�c�YAː    G�b���J��W�疎֗d�T��Ec`?�d��V,9xەP�����g'8ᄹ�5�B^OE?R��+\
��F�����1�F}���L������q�|����c��/�/(xp� H=ch@� 	T���E��eN���B����9,ප(�����(ߏ-Z J�,��@ $%��,@ $�8H;��x�jN�w��m�;��[�;_�.Ӹ_��i%�w��+�Y1�̼]�L���1�4����V��ښj�@m/����C,Vn��y��Bۛ��r&�Z���u&��b/���;_z�n�d+hm�
���,��m�g`"#.���!(�}�D��#i֟ ��<cb�"��M��k�I��1�S�gw;6LO���o7���N��5�js
�Ƒ̚z�&6��*b��[ZZ��Og�򅶵M�>�r�����u2|��	�
$��[<:�e*�a �Ṟ��K�D� �E��H]�$t�BW>ff�B��bӬ���3��[�I�eV*�ǵo�;��ק�_�nA*�g*m^��(���&�W�I͗�b!*@����ZK�f�,Y���O���/�i��σ��p;B�=۟V<b�%j	=i,�!����m���!)�1�STU�6Q\(kϯ�E���aPV�����C��zzkd�H��UX� 6A������~����~��~��G���[���������o���&i7
ؼ��dx@�1l�c��t6W��fR�� �B_W,���Mv�/���qa�Z��B�1I��9[�8zZ�m%3�'R`!�p6F*&�q�
�������ȶ"0�h�C����%Bm� �=���i����ԙ~D4�&�	�D��D�z���G��ၠmD�,w9�-�^q����`o�L����Hѳ�7r���H.���Z�|�6��8&�n]����[���2����e!
�E�a0���<�� 		|"�UW�
ʙ7����L|�Rd�W�! �)FAf����H�E�~�_7��|�7��{�i;p��rB����2�f���	v>�"�!�""��6&�8:���R�%u����$�I$�I$�I$�IxB�K��O�
:�X����*���ߞ��Ol��@gQ
   j
��
"�V�8B���BD!���pl�?������R��]w��M���&�)wh���
z�*+L}��� ��X��6��-ݤXV^ �$Ρ����>��#�;P>�r$x��RW���	3��(�\���� {� �{
E�(�� ���z~l/M�8� H#�R[7��y��K�5V�J/�AH3Dm��I��Gh:뺭�]NС�
|��[���B��u�}� ��:�1p��|��i����r��ߣr�Ԧ�˭e��n���3(�ݏ4� ���-6��w뀧�V&���lW���ۥ�[�_tY��9�'$!ݵ�g]K7���f����ˈ�	��ic09  6�   jP  
�
   ftypjp2     jp2    Ojp2h   ihdr           colr        "cdef                      jp2c�O�Q 2                               �R     �\  PXX`XX`XX`XXXPPX�d  Kakadu-v5.2.1�� 
    5� ������n������gL�)���Ij�:�+g�������(���*hrY����)�96L3*u�%U���,�PY��@��W�����ʦ<�W�^��:����a�(Y��oGV�\��D��;�Ɯ�%���@�L ��{��cO���c`2g��ttO���m�^&s�D(�o��4:�'4~�9�9Ί�I����V�!��\L�A�����o�'撴�;　�½`�Z��FQ/�0�!�M�"~*y��=����v� D p�C��T5ނX�����ed
\]Êf5ωHEr0�~�	��7�N���c��$:�\4��; ������6-űg�W·\U��&��p#N�5G'E:�hx��n¦W��~�`vqbK�2�b��8�\Y������W���Jw������~h �&����F^�誙�)^'Ou�й�1�I���C�[���n��u����b�i����1�k:��+�n8@��?^&}������P�:� �pGq�]>��y>�"b����$��h󌝐�F7k�69B�=����+ᷡvFf�Ǯ�ќ��\�Qbh�'�+�����qso��>75������-3���Z?R����C�o��E�P�ma�������2;;�𡷽A�M
F���祭z����;=h,��,��$�"�(יFQ+m]�X��������?���θp�L({���=�*ߩ��U'��G�5ʈ�A�t7��#/��Eb�W�n �5%�g�,��I�Ow���V"c�����.Fm8+�++�H���f?�%�f'�^ְ�C��Q���ʜ�q�`A�꾪���%JW����<��/a=�ںt���qY�cE�~�P��t���΃" zH#�P@�c鬒��t�"�u� ��;�n�J	T��f�۞b����TRA�
Sȼh����r����	AZ��9���E�t�3N ]~&`_kS��lN���o3Y�/�Sy�~��]P�i{;�/���]�ˉ�J��֟!�a�$��uX�޹r�TK��Kv^0��|��n�tB�E���t�b�X!��l+�<|�ǹ�Ƹr/��>��s_V:�d�SR�R���'�����a�O�^<���V�G�Ȇr1�-�D.෽ք��.R/"S8B�%�(���tID�▣@�ApZ1R�����ےI$�A�<�����J�[Drg�A�$�H��Y�BM�%���������Gk2I$�I&�q{P����2����9��E6�z�;�f��nI$��q!��Hfd7�9Xx��]m�M�^shqy���7$�I$�������([5�TemKw
�x�NR��wxz��N�a�7�&�/�$��(��Gâ@1�����wҏ��^f����n��U�S����uE���4C���P�IٴS'^������g{���|���� p��R�Fw�c�'�Q�Яߓ�>`Z���(�������D?p¶�q������w� /vZ��{�&>@�7)WTa���5��+W K����G��p����.���X�����0�)@��-x1Ł)}�	�]dUi����y"
7�o������4�K�]\'[�i��s��WhO��T�"�-=�W�f�C����ٳ�[������Q�N'�q�0�Ux��*H`)�9�,���Cf�^ʿߡ�Q��9[02���ClijO����Ի�	&�  �w`�o�Q
|�,oȵY��
&-����/߉�a�`��*Hs��ChsV4��]�%҄�Ϡx�6�?=��(�n㝡V���u߸w���[�o��w'�ְ̂=���K����9������J$`��7���2�F��<6:b�V��YPD۟�^\�+��"Tb�u�4�: N���Lű6��֭�����U�WQ� ���a�*/R�Q��n�h �b�ENQ�0�R�DȈ�	�����h��$�i���̣i��/T�Q���
��va� .�m�,��!��_=���q��$����;�pJK�V�"�� ����ǵA /�8}H|��<��|� ��		��,�s-�Dr��
k�FV�E��I!Xi��yH��.������pb������_ ����jsz%#t��GK���@��'
�w	��a<�(��^ɝ�*��vBE*�&;�K�vW*QR���'D�(
�4��~f��Ⱥ�Ȅג�<E����C�W�t��rO����(�8�y��o9�6lZpw��r���O1?�:��?��R�'ɫ�o��X�Ҫ�Zp҇a���E����$��;`����RC��f-gO�0&?ا0~>�����x�tw�P԰Ϧy&������x   E��A߮�O�h'��w�%y�z���&,W�R��O��C��5�k�7�Rµ����g��*Į4|��l��D $ �2]xAyy��:`a��      y� �AC�+c#��5�8jy袻���   Gb̦��HqF�v*Z�����1�Ɩ�Qa�z��K���z�~��)p�{�;#� ����sp��U���|#��o��������q�wSPj��eV�W��"9I߲O="�ͣ�_�&���=®����RM�JMp���fo�f:U#B�1�^����C�?���@��X�d~��N�kl��l@��4�٧����{C���K<�Q|"�7M�[Z:��4�֪N�W��S�}�#���}�bI4cj m�Wwe�K�Z��m��C��s����K�;�%��B��BPERSf���L
��`��,\�VL>��R"��~�m0�/��g�
-�������?��I���x��Ӫ����O`�O2�r��ZEF��.���y0A� 29-eL���V�֘��!�S~x2��#y!�;�$��D�n�'��2jB�Z�ŀ��"f�$_�{���t�b���_P���ʰ���4����{[DU�t$L�G���~gOk����l��bC�a�
��\��;%���Z�6_ଲ��P�+H}��S[@Wp�}�Oήm�̟�/y�� �-m�/�:W�I��Z  ���V����F��  �%m�?�C��+�`9qzG�����nb�B�  tw�$L�?�J��{�:�$`��t����<�8��\�tw��?B���Jf���JKC�k�`�eo����w?�˨�����!��Q��y*�qe�'\�r��,E��Е��R�(�<��W>x�А~	S� k���������O�	v�D�y�,Œ5n�ؐVNY��h S��V/:�y'Ye�r�3�>c��b$Ix�}����]�XN�G���R����{T1�����U�K�4 �0y��=��aG����#pⴶ�5�_��B���  )r2_X��9�K�Vp�P      :�A}�����^o�^�-��4��H�H�T�x�R�dO�l���=/kYi+�:E�B'�C�˸n�Ur�A������0b�8a[��Q1[�� �LZ��Rë��E��?����� �>/�;�ty}�W�(qӱ��7�S�ϩ� �ޖ��fn�!X?
ۯ����o����o���v|ŷV�c���m�vj��S�72;�Q�-Ф )���fv�,4�����]Y�k��`���N��`����f-���V��w~�G��������(8���vC��ݵN���%��ѱ��y��N�J���՛�E���)��r�iQ ��n�x*Rf� ch�[Ň��ȃ	�������|q���G
�T?����X'�Ήpق�_�U��Az��!����̷���kNj��z�~�_7�~n~�%M�u.�P��C�;w�G8��O��i�����1�9D�L�����e�����)r�{��ɾd@�d��/l��N^�Ej9*��l��^��dM\�·�f�d���K�=�2ȸ��ֆx�o����_�����X�;�@|\���ҁ��wf]��֯�t���&(�MՇ1lfߓ�U�-����H5��ZF2��;�V�a����5� �ͧ�@��X�ݒ������2#up�� �G�4���vk`�FK7$@��>�J������b� �m������X�����Y�2z����W�v^]��"�R���Cޮꢝ�&�,�!jx�/���D���e/����J�3�jU��kt�6�����g�4�n���teא�
��@�ٚ�,�	�T\6\U��c�+9����Efo�uFfA�(�W@��!'3i�\zO�/��1㧀�̕�E��Ū����f��P�G��\x�"M�|e�q��6�o�ݰ7-����9�o�E��bd�f����>j-U�>`���a�<6��0Z	�G(�x��h�gn]����[S�����&��3�b:�a,1ku�|�7��|�7��|�Pn�$�=,k�-�f!��1C�`a,YRqF�����/)yK�^R�5���y����+�R򗔼�����K�~�_5�x��c)yK�^R�6���uI�$q��Qo���f'�ku�|ܼ8�B��i�l�'�`X�4-tc�  4��R&�z���^S8�j��'�h�2�T`�F)yL�z�BX��s(����~�$�8�|Qwc��o���M�� �ޤ�� Ҙ�C HKu�HK������V�A�f�wF�����$�`��U���GX�4�ao٨�D����iҖ�Ư�c�b.���{�s��/����+��A-��<�n%=�}[��)����*W{�Z�|�Wm��o�T�WQ|v�@�6�Vl��C�]Lc�2ieiy�{��E�NQ�é�����nb�y�Y�n쐋a���Ʋ��N�
w�[���oA��يLO S,�۵J�ЊN�_�Tޱ~i��@�5y|����=1H��ɡ)���u��򘪪2����C��x�.eY�k���X���Nt�͡O�5�8by�h-�ϐ��[ֆ����U�+[��=�}K�3I����\E�B+z"3�,�A��t���5H����u3mdy�P���� �#�[����, ��?&-8����;�v˷D�b�	6�i�1�v+�F�Q�Χ�:��?�$���2<hAK��W�S������/4�O�{j9�O�an0�峷AQ�k��-�9n�b'����}e1��&OĄ7% >!N���W��؁��Ө��`�G�a�G�����`\ۊrp1���~�ߙ�dRU��X�h���Ev�ۨ�MLG&�&�E�<t!�{ȥ/Q%�����tSD�����ȼf��[���W�`�eº?��;d{���m�C@�y	�%�N� 0����A��R  0�P?M�i����HKk�=�����z�h�>D<�|x���� ��ޱ����  a ��Ybu>H�I $��g�F��A�i����b����-�ALl�D8�X+�:�m�����a�^��]0K��S(��^�bE�B&W|�I֬�!/��М{�z�/$�Z�6xKm�B������b���f�	i��š�}�F�ܺ�V+v��kT�Naiz��>��B�R�K��}1-�_���[�+��pz�/�3�o,Yt.&(�ŢMk�ºz��H�������!9�M��
��Q�t�lV9W�4�P#6-:���nV%����A���*��v|��@�i�Hzȹ��l��qc1���T�`��C�FK2*��t�+ɭ+�w��Ղ���'��r:�iVo��j�7����h�����S�>ėu.Qc��^�h�0�[3�h{�? 4�	��s��"���y��\�S^�a�\%f����1��LZ�6��zB|O�w��V;��YV ��w!ɤz�&;AiH��,�X�����熝��.wҜ���2_"lFT�٥m�r\�΄OIy��G�K�{.�9ݍ�`�v��;š�~�W�D�I.�U���Z�n#�_qf}��"+���Hr8�g��R���8�[dY<G�."�
J�in�S��������径 un������"��o�#��kҙW�9���W�L��9� �*����J>q�J�d�ra�
>�E����P�m��R?j������Zo�Nq>���JO�B}B�o���%�Twu4�ӆ�9@�a!�+�:��0;-`�+n�o����o����o��CM�XE��U˼~T	(����AS|�f�|�.H�:, i�[�?ExYg"z*Ҕ�8AՂW����@\:��P  ��薷�>��P�$�ڲISă���j�a)�	�Y�44m��O�m���j�L�y:X�\1Xd���GN��?��>%^3�&Ƹ�Hj�$܊+�0�-͎� �$IG���f�Ћ���-��:4�t�K�7���������n]����[P�U}��Mv 0�����\g�O��Иb�����o����o��gI'V}_L��, ��l`荗X���/��7������i}87�HIh�/��� ������o����o��bPX�>ځ���.*	���=R��+n�o����o����E�rB���u������ H8W��H�_��� �B_b�}Ϗ<�{��d�      �xB���?X8i�GB�9���w�k0ٹ��E%w�ś�+0�   � ~G���jy�����֩0§�{K�	�cI�eyB� ���.nkm}t���A�j�'��"��%��?��_F\��i�ED�E�`��#��~��g/�Y���?��<O���>��#�;D@#�|Ca�	*��ȭ2�?����ZQ_[�A����� $�1x9o�� ��s�-/$M	��� $f}�x ��C�/d�/�P�o���ۀ a {�� �mⓖ�o�Gw;"��Y�Х蛘�כ6Kڿ�dīȂ�Ġ^��^�1�W�
���KS�ip6�(����܁�@`9��XPJKSE��8�ߖj0�gH�w]�����j�p?b��FLO��K�[�_�-��D�S��/Z�\oH�0�OQ���bcЌ��Lb�:۾&�k+�9ߠ�o}�8�3�
���՘�����x1R!Ӟ`��x�������u��4����w�����i:�?�?��/�?�G�p��ud
��i�X�do[h���A�?�ۉ��_��O�hq�{�*yP*��~�p�6*���ZD��axD�b�����o����o���E5�+n�o��վ��"1=`�[�����s� �b�~�)ҥ��q���t���(N��\`Hp�I5��S��<l���oVVq��3}�)(P�FH���9����So��I�W8=��z�vN���7Ubo�Mw���8H��s����F����Z�H�t���#��n:X+�9��Z�I��(ұmպ�+/�D*d(^����H��&���s��������1oJ+�I�f%ٌfض��Ծ�\J��&�����D�T����V`����&�.��jm��E�Ll8E��$��r�>�̲W���>����u���Ga��<�A�f��\�AVR��^��]��]M ��ڃ}LX��:��&3�%T8�GOF�UabA���<�}p����5��t�p�ͦ�?s)L��J��7��@8I�	Q=��$��+�p���|f�*�.��J�|��
�z4
Ģ�y��t�+�R��A�Ҧ*iM0���oLb9�;���V/��*s^�!Zh��GՠY��Z�Sy�<�w��a�xĈ��:1�+kٵ\ y�19֟�3G�P�)>u��fn�Xyqt,�P�>o��tK1:[�,�DZ�T�.B���nYb�_��ᚲ��Z��撻��q�YQ���],"�LZt�bN�_��#�Ev)��t`5R<ӽ �.Ô��3�Y���`%�:88�2�OK��X���m��|(���L�χѺ��8o���D�_��{��Sr�����DF�? Jx���Z���ʥ[u��=��5�׀<�<^�o������/t�|�a�y�̰���Y7p�;��*V�"���?��	��'�[�kG��J���]�X4��A$W�j��^�qi5�;Lx��q47���E����<+��eu�� D0�@X%Z�WF�u@� =�S��p� �u!Z2D�$���#���V,}�JJ0�l�#�,`�t����gi���&�w��a共=����K�Kᖬ:XwXU�U�,��o+��f!j�P����hD �Ƴ�<������>*��d�� ��lS1֋$�7E��M����%(�z\P&n�K:i�5p�����x,��Т�,�[u�|�7�2
�a�[��	k���n���剂���=�p���K$���٭.BO��|�ߕlUa��6�}l��`��G;M����-�U��ּ�5�<��E����΄ٵ+U�Q��#���c#N@N���/��K��̀���V��������i��:��M՘����+�Q0=0��d5��B�#W���6'�9lt6��q���(�(,d> �j�d?愉"�9j&QJ6��se��&i�Z�|�7��|�7�zk�1n;�J3�Ҟ�m���|�7˃Y��ރ�x<P{UH���DՂ�s�q	��+n�o�7�X�QQ�	�D����3W"�oq��řPCب7QQtyS�O}HE���K.�E�$�sHR�!h���VD{[��R��d�����T�D�|`oU���!��x�q��/0��1͎���rJᢖ�5p������ ��u���E����j�,)�"�~�݌q���(�޳�czGa�P���o����o����o�R��7��|�7��|�7��|�7﫮�o����o����o����o����V�|�7��Y~iZ�HNܰŭ��H���<�H��5��@Bڎf��s��es�l�h4��0��4�NF��Q.:��E���gM�����������`���-� �	�~�| �� 		~� HH��E?��󖌐lW�ld#q���&���MA������?2���*d��F��>�߆w�RAyUI-t��J>�=��R$�S���S�Ώ����L��x�ٳv�@7�F9<���2U8�������"�
[���ۅ�L�
{$�j���f�ii�����-��ȕ'��O����rC�ڕ�y��w��8(��IO��*DJ=+ES�8	��vq5<���l�	��
��_M���np�S<�lH�=���+ ���}��4#eՖ���5~0��*{BQ�$��A����p�j��i-�D���U3��4��RO��p��/i� !�jP�l�V[b�=�X�4�4�j4�zT��Ӏ�$�y[n�-�]|��s;���a!raz\�bpy!%[��?+��O(��~�)+=l�f=�Ff�#�!Л:`ɡ|��j����EtiP�w��1�ןr}�&�d���Nn�#�mkɰ0���x�M�����O�#�f� ���USf0��~2�ڂQt����E���IB�� �����^2�+fn
y�7$hk"|��z?��7犇�?�(�~{�V����4�yJ���J��5jXľ�4�Ņ�{�Մ��I��H�!"}��qxL�!彔)�*3~�f՗�m;��9d2��	Y�c����^:������L�ON�8�o��QK��
�lt����?P�t=4����o�%=_5�YR.u����'�� ���$=>~��]a�ZXh�*u��/���֠���;oO
 J;v��ڌ���$���Ɂ�pb���簙I�߮X�$[�M��Ѣ��_)i��c(~�X��G����3`������F���P�[��؁� �J�~�t'!|��y���؋� \DhD��0�%�,2�L����m��}o6c�0�k;�<��:S��v�r�K�w��|A�B�0�$��/F�U��Nr&?|�U6~�]���÷�V^����(3zLA��6q���l�2�ˏ�:U��76)��瀒���1�l-x�(n�z>%�����6�MV��ސ*�0����!�Q귗<d��	4_�B�����V)y�_��d�IW��N-%*�G����)�آX��9Z�����^�i�f��"I,@�S�ǿ����Q�����Sk!u��b���Hw2��X Y����A�84�d#�y- ���g����TCN��KWvJBdo�B0�����o�+��(��{�I^��~����~��G�c�����-�֓;�\ɠ�,ف�G��.�rȶ,�2����P��#r���)y��v�G���s��u58���`��ԡ�ei��v[��ܹvIFȶeK�e8-�����h��c6د3&8RM̙Nn`��S����)@��P���`'�GU<���EL(���lliN��}>�a*�с�6��>�J������Z>K���>��"aG�

B�>��"aG�

B�>��l|�G��Rh��[�Q𩳶L��B���n��_ �I�(#�[$�(#�S�m��)����)��� �:#f���t  HK���  		GE����ģ		 �BOqc		 �BNWc		 �BF�� �:#f���t  HK���  		GE����ģ		 �BOqc		 �BNWc		 �BF�� �^�x����D�$m��  #ȁ�c�U�_H����W���?xVLw�a���
���-WV��q���>����J��>q�H�ʆ.���L�_쩤	�(��
^M��#W9�|o��M��>I�ķ�d\S]�&�(D��f���2� ؟�]�Y۫<���X��޳o�^�\��q(�;�N�	%G��}w���zj^<MdͮV�u�[�p�+��}�b�I�V�������2c���m���V�SIl��)�dSU�{�rYU�$����cb_m!#\r�Ct����1S5�6�" ��p��(���<���P���-.8�5��;�Y��q�>�q?�,0 �+�u���|���	�& {��jӖ�
�V�f �5^J��.���L��!�2�.���d�x���t�?����Pvif�j�MI��](�x:�2�\�!B�!TEA��P���]�A�,�E����Q:M�Kp!rNhO� ���){!��/��X!I�w�ߺ�2�4{���QP���'�̖en�5�f�Ԣ��X�U�Ӹ[;��dhM�e^;`k�	d�����ቼ�X-��Ɣ��ՠA����u߅�#��R����c����k*ñ�9>��z���`5�r;��8��0��c
&$\J;����գ�����y�d��a	�"�)>�����\B������@��B�T⛍����4j)��>�������.W�y�7��	��7�������+fֻ�p[�)�z7L���ф�j*�"/�TD9#.{����L׶pv���y���<<|��Akp����>��&��g5S����Z��u>�ɖ�����I5C�����_��5�A��}s���z�y��h	PЂ߇��Y �.�gμ5��'�<�B�1�����4�(b���YR������Pj�T�?k�>��V� �|Hu�ÍUR=�+���v���بo$*���rcJ��>�U0�I�#&�� �^c�ڄ��m��r-^�槶�Y-
|T+j��~[rx2�!����+����knR48�� Klw�b�K�?,�p�͕��O�$?�q^T*��]�ә���9��3����a��_��%z�Ri���AD��������8@�'��'�9)q�Ɗ�K����z����X���ďQ~�_�����i3�t�/g�j��矐�Jy�h��$p���Xj�,�)B�q5��'��i�
��ܽ�y�k��(B����}��ag!�%��a���j�llR��EB��~����`C�����I 䡡�I�/���.��] ;W����Z��g�vYmg+���9'��1�H�!�t��"n��� � �]̪ � 8��]��T=�4�����|���G��'�j�4eiw�C?jo�a�E�m�/�\_Qt��y�G�w��p�P�����a��K���!�t+`�0@�~P���xэ���M�D�=��� 6�)F�8��3_�jC�5�����A��s%��m����l�95�/Z=�#8i�;��#�?��o�T��x =���T�+v�P�(�L���c2{�u:�NR��@i��a��~� L]I�k�=�bJ�8��
�sF�����gD�o�ca�x��� .9a+���z)����L	@�f���#Dg�Ko^�h�x*�������h>;	��ĵ/��1O�,gpe��h �E�ň�ٮ�yn���P���/�/��ɨ�eP�s� ������W�Ǌr�T��$���X���ӳV�&�|��]}��Y��y��4mTQ��l6��a��l5��	Dp�,��1O�,gpe��h �E�ň�ٮ���1��.��  �BBL��bHK���0��I�-n�o����o����o���1O���)aK�q�$d!J�����Z��L�&�	��Y�HK&3gBێE�U�=d4�I�D��E������1���R��������mnU�XH:�h�%-q��9�-X ��[j�^��J��L��'��a`?
ۯ����o���9N��E�����a��6����qV{� c�ެR;��+6z����.�
� �	�~����� $$��"1��� ��9X�0����R�
���{��N���~�x/`B�-A�|y�ò�͈P���}7p��{�̺cK����D�P����%�sP��fei���a�Ɔ�����n��|��w�����yhn)	�i<��Rz]~���17���o������qtL�z��S-�l�#h�	j�� iv�n��n���^S��d�u�h3C[�1��>8�c}�ie�2��r��WL� �]�e�H#B����ƗS�{�v�������j1�kPح�K�K�0��GOv��~�'�}�\5�5�~[�al�+�}'
	AP����"F���{�����M`��1����及s��;`���B٩�l 0�0?���eX���2vݰ�E�� ~Ç��� �:#�.@ $%�HJ$������� �:#�.@ $%�HJ$������� �^�u��ղH"�-�<ʝm��s��g�H�0�b��+"a��K5�r:�`��=[������
RY�$4JKʗ1����aO��5�/�o����Q��J�R���<0��;U]�2�a�Hڃ��w|(2�|�A��4��\�ؤ�     ��Uj�2���)���r-"�D�v�S�X��=�َ�� � Eǅc88^[ƹg�a���Ѷ�6^�]`k�KS�c����hd�6I�h������.���7�a�^�l�*��u#3,]���
U ��� 1J+���JV��־��s�s4Tr5�6�/jS��[x�ɐ�Ma��������8�}��/d�xI)JL�o�SYrY@��{~�乙!B&�dh�>�훸Ot&�H�"%�ҷ�]��2/�S����ѓ�""n-H�LhwIBx�^Xa�%�|4��D
p�fX��$���$0�_�ٲ���O�� �        �   Macintosh HD               �{�H+   ���
hfr.nc.cdl                                                      ��'�ic?        ����  	                	test_data     �{<�      �i��      ��� ��q ��� +ȳ +Ǫ 	� �S :�  \Macintosh HD:Users:cmueller:Development:OOI:Dev:datamodel:pytaps-ptypes:test_data:hfr.nc.cdl   
 h f r . n c . c d l    M a c i n t o s h   H D  OUsers/cmueller/Development/OOI/Dev/datamodel/pytaps-ptypes/test_data/hfr.nc.cdl   /    ��  �   ����            �         `        �         D         �         �         �         �          $      0   P      �  �      �         �  �      �  X      �  �        �  d       �  p�      