netcdf roms {
dimensions:
	ocean_time = 3 ;
	s_w = 37 ;
	eta_rho = 82 ;
	xi_rho = 130 ;
	tracer = 2 ;
	s_rho = 36 ;
	eta_u = 82 ;
	xi_u = 129 ;
	eta_v = 81 ;
	xi_v = 130 ;
	boundary = 4 ;
	eta_psi = 81 ;
	xi_psi = 129 ;
	maxStrlen64 = 64 ;
variables:
	float AKs(ocean_time, s_w, eta_rho, xi_rho) ;
		AKs:long_name = "time-averaged salinity vertical diffusion coefficient" ;
		AKs:units = "meter2 second-1" ;
		AKs:time = "ocean_time" ;
		AKs:coordinates = "lon_rho lat_rho s_w ocean_time" ;
		AKs:field = "AKs, scalar, series" ;
		AKs:_FillValue = 1.e+37f ;
	float AKt(ocean_time, s_w, eta_rho, xi_rho) ;
		AKt:long_name = "time-averaged temperature vertical diffusion coefficient" ;
		AKt:units = "meter2 second-1" ;
		AKt:time = "ocean_time" ;
		AKt:coordinates = "lon_rho lat_rho s_w ocean_time" ;
		AKt:field = "AKt, scalar, series" ;
		AKt:_FillValue = 1.e+37f ;
	float AKv(ocean_time, s_w, eta_rho, xi_rho) ;
		AKv:long_name = "time-averaged vertical viscosity coefficient" ;
		AKv:units = "meter2 second-1" ;
		AKv:time = "ocean_time" ;
		AKv:coordinates = "lon_rho lat_rho s_w ocean_time" ;
		AKv:field = "AKv, scalar, series" ;
		AKv:_FillValue = 1.e+37f ;
	double Akk_bak ;
		Akk_bak:long_name = "background vertical mixing coefficient for turbulent energy" ;
		Akk_bak:units = "meter2 second-1" ;
	double Akp_bak ;
		Akp_bak:long_name = "background vertical mixing coefficient for length scale" ;
		Akp_bak:units = "meter2 second-1" ;
	double Akt_bak(tracer) ;
		Akt_bak:long_name = "background vertical mixing coefficient for tracers" ;
		Akt_bak:units = "meter2 second-1" ;
	double Akv_bak ;
		Akv_bak:long_name = "background vertical mixing coefficient for momentum" ;
		Akv_bak:units = "meter2 second-1" ;
	double Charnok_alpha ;
		Charnok_alpha:long_name = "Charnok factor for surface roughness" ;
	double CrgBan_cw ;
		CrgBan_cw:long_name = "surface flux due to Craig and Banner wave breaking" ;
	double Cs_r(s_rho) ;
		Cs_r:long_name = "S-coordinate stretching curves at RHO-points" ;
		Cs_r:valid_min = -1. ;
		Cs_r:valid_max = 0. ;
		Cs_r:field = "Cs_r, scalar" ;
	double Cs_w(s_w) ;
		Cs_w:long_name = "S-coordinate stretching curves at W-points" ;
		Cs_w:valid_min = -1. ;
		Cs_w:valid_max = 0. ;
		Cs_w:field = "Cs_w, scalar" ;
	float DU_avg1(ocean_time, eta_u, xi_u) ;
		DU_avg1:long_name = "time averaged u-flux for 2D equations" ;
		DU_avg1:units = "meter3 second-1" ;
		DU_avg1:time = "ocean_time" ;
		DU_avg1:coordinates = "lon_u lat_u ocean_time" ;
		DU_avg1:field = "DU_avg1, scalar, series" ;
		DU_avg1:_FillValue = 1.e+37f ;
	float DU_avg2(ocean_time, eta_u, xi_u) ;
		DU_avg2:long_name = "time averaged u-flux for 3D equations coupling" ;
		DU_avg2:units = "meter3 second-1" ;
		DU_avg2:time = "ocean_time" ;
		DU_avg2:coordinates = "lon_u lat_u ocean_time" ;
		DU_avg2:field = "DU_avg2, scalar, series" ;
		DU_avg2:_FillValue = 1.e+37f ;
	float DV_avg1(ocean_time, eta_v, xi_v) ;
		DV_avg1:long_name = "time averaged v-flux for 2D equations" ;
		DV_avg1:units = "meter3 second-1" ;
		DV_avg1:time = "ocean_time" ;
		DV_avg1:coordinates = "lon_v lat_v ocean_time" ;
		DV_avg1:field = "DV_avg1, scalar, series" ;
		DV_avg1:_FillValue = 1.e+37f ;
	float DV_avg2(ocean_time, eta_v, xi_v) ;
		DV_avg2:long_name = "time averaged v-flux for 3D equations coupling" ;
		DV_avg2:units = "meter3 second-1" ;
		DV_avg2:time = "ocean_time" ;
		DV_avg2:coordinates = "lon_v lat_v ocean_time" ;
		DV_avg2:field = "DV_avg2, scalar, series" ;
		DV_avg2:_FillValue = 1.e+37f ;
	double FSobc_in(boundary) ;
		FSobc_in:long_name = "free-surface inflow, nudging inverse time scale" ;
		FSobc_in:units = "second-1" ;
	double FSobc_out(boundary) ;
		FSobc_out:long_name = "free-surface outflow, nudging inverse time scale" ;
		FSobc_out:units = "second-1" ;
	double Falpha ;
		Falpha:long_name = "Power-law shape barotropic filter parameter" ;
	double Fbeta ;
		Fbeta:long_name = "Power-law shape barotropic filter parameter" ;
	double Fgamma ;
		Fgamma:long_name = "Power-law shape barotropic filter parameter" ;
	int LtracerSrc(tracer) ;
		LtracerSrc:long_name = "tracer point sources and simck activation switch" ;
		LtracerSrc:flag_values = 0, 1 ;
		LtracerSrc:flag_meanings = ".FALSE. .TRUE." ;
	double M2nudg ;
		M2nudg:long_name = "2D momentum nudging/relaxation inverse time scale" ;
		M2nudg:units = "day-1" ;
	double M2obc_in(boundary) ;
		M2obc_in:long_name = "2D momentum inflow, nudging inverse time scale" ;
		M2obc_in:units = "second-1" ;
	double M2obc_out(boundary) ;
		M2obc_out:long_name = "2D momentum outflow, nudging inverse time scale" ;
		M2obc_out:units = "second-1" ;
	double M3nudg ;
		M3nudg:long_name = "3D momentum nudging/relaxation inverse time scale" ;
		M3nudg:units = "day-1" ;
	double M3obc_in(boundary) ;
		M3obc_in:long_name = "3D momentum inflow, nudging inverse time scale" ;
		M3obc_in:units = "second-1" ;
	double M3obc_out(boundary) ;
		M3obc_out:long_name = "3D momentum outflow, nudging inverse time scale" ;
		M3obc_out:units = "second-1" ;
	double Tcline ;
		Tcline:long_name = "S-coordinate surface/bottom layer width" ;
		Tcline:units = "meter" ;
	double Tnudg(tracer) ;
		Tnudg:long_name = "Tracers nudging/relaxation inverse time scale" ;
		Tnudg:units = "day-1" ;
	double Tobc_in(boundary, tracer) ;
		Tobc_in:long_name = "tracers inflow, nudging inverse time scale" ;
		Tobc_in:units = "second-1" ;
	double Tobc_out(boundary, tracer) ;
		Tobc_out:long_name = "tracers outflow, nudging inverse time scale" ;
		Tobc_out:units = "second-1" ;
	int Vstretching ;
		Vstretching:long_name = "vertical terrain-following stretching function" ;
	int Vtransform ;
		Vtransform:long_name = "vertical terrain-following transformation equation" ;
	double Znudg ;
		Znudg:long_name = "free-surface nudging/relaxation inverse time scale" ;
		Znudg:units = "day-1" ;
	double Zob ;
		Zob:long_name = "bottom roughness" ;
		Zob:units = "meter" ;
	double Zos ;
		Zos:long_name = "surface roughness" ;
		Zos:units = "meter" ;
	double Zos_hsig_alpha ;
		Zos_hsig_alpha:long_name = "wave amplitude factor for surface roughness" ;
	double angle(eta_rho, xi_rho) ;
		angle:long_name = "angle between XI-axis and EAST" ;
		angle:units = "radians" ;
		angle:coordinates = "lon_rho lat_rho" ;
		angle:field = "angle, scalar" ;
	double dstart ;
		dstart:long_name = "time stamp assigned to model initilization" ;
		dstart:units = "days since 2006-01-01 00:00:00" ;
	double dt ;
		dt:long_name = "size of long time-steps" ;
		dt:units = "second" ;
	double dtfast ;
		dtfast:long_name = "size of short time-steps" ;
		dtfast:units = "second" ;
	double el ;
		el:long_name = "domain length in the ETA-direction" ;
		el:units = "meter" ;
	double f(eta_rho, xi_rho) ;
		f:long_name = "Coriolis parameter at RHO-points" ;
		f:units = "second-1" ;
		f:coordinates = "lon_rho lat_rho" ;
		f:field = "coriolis, scalar" ;
	double gamma2 ;
		gamma2:long_name = "slipperiness parameter" ;
	double gls_Kmin ;
		gls_Kmin:long_name = "minimum value of specific turbulent kinetic energy" ;
	double gls_Pmin ;
		gls_Pmin:long_name = "minimum Value of dissipation" ;
	double gls_c1 ;
		gls_c1:long_name = "shear production coefficient" ;
	double gls_c2 ;
		gls_c2:long_name = "dissipation coefficient" ;
	double gls_c3m ;
		gls_c3m:long_name = "buoyancy production coefficient (minus)" ;
	double gls_c3p ;
		gls_c3p:long_name = "buoyancy production coefficient (plus)" ;
	double gls_cmu0 ;
		gls_cmu0:long_name = "stability coefficient" ;
	double gls_m ;
		gls_m:long_name = "turbulent kinetic energy exponent" ;
	double gls_n ;
		gls_n:long_name = "turbulent length scale exponent" ;
	double gls_p ;
		gls_p:long_name = "stability exponent" ;
	double gls_sigk ;
		gls_sigk:long_name = "constant Schmidt number for TKE" ;
	double gls_sigp ;
		gls_sigp:long_name = "constant Schmidt number for PSI" ;
	double h(eta_rho, xi_rho) ;
		h:long_name = "bathymetry at RHO-points" ;
		h:units = "meter" ;
		h:coordinates = "lon_rho lat_rho" ;
		h:field = "bath, scalar" ;
	double hc ;
		hc:long_name = "S-coordinate parameter, critical depth" ;
		hc:units = "meter" ;
	double lat_psi(eta_psi, xi_psi) ;
		lat_psi:long_name = "latitude of PSI-points" ;
		lat_psi:units = "degree_north" ;
		lat_psi:standard_name = "latitude" ;
		lat_psi:field = "lat_psi, scalar" ;
	double lat_rho(eta_rho, xi_rho) ;
		lat_rho:long_name = "latitude of RHO-points" ;
		lat_rho:units = "degree_north" ;
		lat_rho:standard_name = "latitude" ;
		lat_rho:field = "lat_rho, scalar" ;
	double lat_u(eta_u, xi_u) ;
		lat_u:long_name = "latitude of U-points" ;
		lat_u:units = "degree_north" ;
		lat_u:standard_name = "latitude" ;
		lat_u:field = "lat_u, scalar" ;
	double lat_v(eta_v, xi_v) ;
		lat_v:long_name = "latitude of V-points" ;
		lat_v:units = "degree_north" ;
		lat_v:standard_name = "latitude" ;
		lat_v:field = "lat_v, scalar" ;
	double lon_psi(eta_psi, xi_psi) ;
		lon_psi:long_name = "longitude of PSI-points" ;
		lon_psi:units = "degree_east" ;
		lon_psi:standard_name = "longitude" ;
		lon_psi:field = "lon_psi, scalar" ;
	double lon_rho(eta_rho, xi_rho) ;
		lon_rho:long_name = "longitude of RHO-points" ;
		lon_rho:units = "degree_east" ;
		lon_rho:standard_name = "longitude" ;
		lon_rho:field = "lon_rho, scalar" ;
	double lon_u(eta_u, xi_u) ;
		lon_u:long_name = "longitude of U-points" ;
		lon_u:units = "degree_east" ;
		lon_u:standard_name = "longitude" ;
		lon_u:field = "lon_u, scalar" ;
	double lon_v(eta_v, xi_v) ;
		lon_v:long_name = "longitude of V-points" ;
		lon_v:units = "degree_east" ;
		lon_v:standard_name = "longitude" ;
		lon_v:field = "lon_v, scalar" ;
	double mask_psi(eta_psi, xi_psi) ;
		mask_psi:long_name = "mask on psi-points" ;
		mask_psi:flag_values = 0., 1. ;
		mask_psi:flag_meanings = "land water" ;
		mask_psi:coordinates = "lon_psi lat_psi" ;
	double mask_rho(eta_rho, xi_rho) ;
		mask_rho:long_name = "mask on RHO-points" ;
		mask_rho:flag_values = 0., 1. ;
		mask_rho:flag_meanings = "land water" ;
		mask_rho:coordinates = "lon_rho lat_rho" ;
	double mask_u(eta_u, xi_u) ;
		mask_u:long_name = "mask on U-points" ;
		mask_u:flag_values = 0., 1. ;
		mask_u:flag_meanings = "land water" ;
		mask_u:coordinates = "lon_u lat_u" ;
	double mask_v(eta_v, xi_v) ;
		mask_v:long_name = "mask on V-points" ;
		mask_v:flag_values = 0., 1. ;
		mask_v:flag_meanings = "land water" ;
		mask_v:coordinates = "lon_v lat_v" ;
	int nAVG ;
		nAVG:long_name = "number of time-steps between time-averaged records" ;
	int nHIS ;
		nHIS:long_name = "number of time-steps between history records" ;
	int nRST ;
		nRST:long_name = "number of time-steps between restart records" ;
	int ndefAVG ;
		ndefAVG:long_name = "number of time-steps between the creation of average files" ;
	int ndefHIS ;
		ndefHIS:long_name = "number of time-steps between the creation of history files" ;
	int ndtfast ;
		ndtfast:long_name = "number of short time-steps" ;
	double nl_tnu2(tracer) ;
		nl_tnu2:long_name = "nonlinear model Laplacian mixing coefficient for tracers" ;
		nl_tnu2:units = "meter2 second-1" ;
	double nl_visc2 ;
		nl_visc2:long_name = "nonlinear model Laplacian mixing coefficient for momentum" ;
		nl_visc2:units = "meter2 second-1" ;
	int ntimes ;
		ntimes:long_name = "number of long time-steps" ;
	int ntsAVG ;
		ntsAVG:long_name = "starting time-step for accumulation of time-averaged fields" ;
	double ocean_time(ocean_time) ;
		ocean_time:long_name = "averaged time since initialization" ;
		ocean_time:units = "seconds since 2006-01-01 00:00:00" ;
		ocean_time:calendar = "gregorian" ;
		ocean_time:field = "time, scalar, series" ;
	double pm(eta_rho, xi_rho) ;
		pm:long_name = "curvilinear coordinate metric in XI" ;
		pm:units = "meter-1" ;
		pm:coordinates = "lon_rho lat_rho" ;
		pm:field = "pm, scalar" ;
	double pn(eta_rho, xi_rho) ;
		pn:long_name = "curvilinear coordinate metric in ETA" ;
		pn:units = "meter-1" ;
		pn:coordinates = "lon_rho lat_rho" ;
		pn:field = "pn, scalar" ;
	double rdrg ;
		rdrg:long_name = "linear drag coefficient" ;
		rdrg:units = "meter second-1" ;
	double rdrg2 ;
		rdrg2:long_name = "quadratic drag coefficient" ;
	double rho0 ;
		rho0:long_name = "mean density used in Boussinesq approximation" ;
		rho0:units = "kilogram meter-3" ;
	double s_rho(s_rho) ;
		s_rho:long_name = "S-coordinate at RHO-points" ;
		s_rho:valid_min = -1. ;
		s_rho:valid_max = 0. ;
		s_rho:positive = "up" ;
		s_rho:standard_name = "ocean_s_coordinate_g1" ;
		s_rho:formula_terms = "s: s_rho C: Cs_r eta: zeta depth: h depth_c: hc" ;
		s_rho:field = "s_rho, scalar" ;
	double s_w(s_w) ;
		s_w:long_name = "S-coordinate at W-points" ;
		s_w:valid_min = -1. ;
		s_w:valid_max = 0. ;
		s_w:positive = "up" ;
		s_w:standard_name = "ocean_s_coordinate_g1" ;
		s_w:formula_terms = "s: s_w C: Cs_w eta: zeta depth: h depth_c: hc" ;
		s_w:field = "s_w, scalar" ;
	float salt(ocean_time, s_rho, eta_rho, xi_rho) ;
		salt:long_name = "time-averaged salinity" ;
		salt:time = "ocean_time" ;
		salt:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		salt:field = "salinity, scalar, series" ;
		salt:_FillValue = 1.e+37f ;
	float shflux(ocean_time, eta_rho, xi_rho) ;
		shflux:long_name = "time-averaged surface net heat flux" ;
		shflux:units = "watt meter-2" ;
		shflux:negative_value = "upward flux, cooling" ;
		shflux:positive_value = "downward flux, heating" ;
		shflux:time = "ocean_time" ;
		shflux:coordinates = "lon_rho lat_rho ocean_time" ;
		shflux:field = "surface heat flux, scalar, series" ;
		shflux:_FillValue = 1.e+37f ;
	char spherical(maxStrlen64) ;
		spherical:long_name = "grid type logical switch" ;
		spherical:flag_values = "T, F" ;
		spherical:flag_meanings = "spherical Cartesian" ;
	float sustr(ocean_time, eta_u, xi_u) ;
		sustr:long_name = "time-averaged surface u-momentum stress" ;
		sustr:units = "newton meter-2" ;
		sustr:time = "ocean_time" ;
		sustr:coordinates = "lon_u lat_u ocean_time" ;
		sustr:field = "surface u-momentum stress, scalar, series" ;
		sustr:_FillValue = 1.e+37f ;
	float svstr(ocean_time, eta_v, xi_v) ;
		svstr:long_name = "time-averaged surface v-momentum stress" ;
		svstr:units = "newton meter-2" ;
		svstr:time = "ocean_time" ;
		svstr:coordinates = "lon_v lat_v ocean_time" ;
		svstr:field = "surface v-momentum stress, scalar, series" ;
		svstr:_FillValue = 1.e+37f ;
	float swrad(ocean_time, eta_rho, xi_rho) ;
		swrad:long_name = "time-averaged solar shortwave radiation flux" ;
		swrad:units = "watt meter-2" ;
		swrad:negative_value = "upward flux, cooling" ;
		swrad:positive_value = "downward flux, heating" ;
		swrad:time = "ocean_time" ;
		swrad:coordinates = "lon_rho lat_rho ocean_time" ;
		swrad:field = "shortwave radiation, scalar, series" ;
		swrad:_FillValue = 1.e+37f ;
	double sz_alpha ;
		sz_alpha:long_name = "surface flux from wave dissipation" ;
	float temp(ocean_time, s_rho, eta_rho, xi_rho) ;
		temp:long_name = "time-averaged potential temperature" ;
		temp:units = "Celsius" ;
		temp:time = "ocean_time" ;
		temp:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		temp:field = "temperature, scalar, series" ;
		temp:_FillValue = 1.e+37f ;
	double theta_b ;
		theta_b:long_name = "S-coordinate bottom control parameter" ;
	double theta_s ;
		theta_s:long_name = "S-coordinate surface control parameter" ;
	float u(ocean_time, s_rho, eta_u, xi_u) ;
		u:long_name = "time-averaged u-momentum component" ;
		u:units = "meter second-1" ;
		u:time = "ocean_time" ;
		u:coordinates = "lon_u lat_u s_rho ocean_time" ;
		u:field = "u-velocity, scalar, series" ;
		u:_FillValue = 1.e+37f ;
	float ubar(ocean_time, eta_u, xi_u) ;
		ubar:long_name = "time-averaged vertically integrated u-momentum component" ;
		ubar:units = "meter second-1" ;
		ubar:time = "ocean_time" ;
		ubar:coordinates = "lon_u lat_u ocean_time" ;
		ubar:field = "ubar-velocity, scalar, series" ;
		ubar:_FillValue = 1.e+37f ;
	float v(ocean_time, s_rho, eta_v, xi_v) ;
		v:long_name = "time-averaged v-momentum component" ;
		v:units = "meter second-1" ;
		v:time = "ocean_time" ;
		v:coordinates = "lon_v lat_v s_rho ocean_time" ;
		v:field = "v-velocity, scalar, series" ;
		v:_FillValue = 1.e+37f ;
	float vbar(ocean_time, eta_v, xi_v) ;
		vbar:long_name = "time-averaged vertically integrated v-momentum component" ;
		vbar:units = "meter second-1" ;
		vbar:time = "ocean_time" ;
		vbar:coordinates = "lon_v lat_v ocean_time" ;
		vbar:field = "vbar-velocity, scalar, series" ;
		vbar:_FillValue = 1.e+37f ;
	float w(ocean_time, s_w, eta_rho, xi_rho) ;
		w:long_name = "time-averaged vertical momentum component" ;
		w:units = "meter second-1" ;
		w:time = "ocean_time" ;
		w:coordinates = "lon_rho lat_rho s_w ocean_time" ;
		w:field = "w-velocity, scalar, series" ;
		w:_FillValue = 1.e+37f ;
	double xl ;
		xl:long_name = "domain length in the XI-direction" ;
		xl:units = "meter" ;
	float zeta(ocean_time, eta_rho, xi_rho) ;
		zeta:long_name = "time-averaged free-surface" ;
		zeta:units = "meter" ;
		zeta:time = "ocean_time" ;
		zeta:coordinates = "lon_rho lat_rho ocean_time" ;
		zeta:field = "free-surface, scalar, series" ;
		zeta:_FillValue = 1.e+37f ;

// global attributes:
		:file = "espresso_avg_2254_0006.nc" ;
		:format = "netCDF-3 classic file" ;
		:Conventions = "CF-1.0" ;
		:type = "ROMS/TOMS averages file" ;
		:title = "ESPRESSO" ;
		:rst_file = "espresso_rst_2254.nc" ;
		:his_base = "espresso_his_2254" ;
		:avg_base = "espresso_avg_2254" ;
		:grd_file = "/home/om/roms/espresso/Data/espresso_grid_c05.nc" ;
		:ini_file = "/home/julia/ROMS/espresso/RealTime/Storage/run03/espresso_ini_2254.nc" ;
		:frc_file_01 = "/home/om/roms/espresso/Data/espresso_tide_c05_20060101.nc" ;
		:frc_file_02 = "../Data/espresso_river_20030101_now.nc" ;
		:frc_file_03 = "../Data/rain_ncepnam_3hourly_MAB_and_GoM.nc" ;
		:frc_file_04 = "../Data/swrad_ncepnam_3hourly_MAB_and_GoM.nc" ;
		:frc_file_05 = "../Data/Tair_ncepnam_3hourly_MAB_and_GoM.nc" ;
		:frc_file_06 = "../Data/Pair_ncepnam_3hourly_MAB_and_GoM.nc" ;
		:frc_file_07 = "../Data/Qair_ncepnam_3hourly_MAB_and_GoM.nc" ;
		:frc_file_08 = "../Data/lwrad_ncepnam_3hourly_MAB_and_GoM.nc" ;
		:frc_file_09 = "../Data/Uwind_ncepnam_3hourly_MAB_and_GoM.nc" ;
		:frc_file_10 = "../Data/Vwind_ncepnam_3hourly_MAB_and_GoM.nc" ;
		:bry_file = "../Data/espresso_bdry.nc" ;
		:clm_file = "../Data/espresso_clm.nc" ;
		:script_file = "nl_ocean_espresso.in" ;
		:svn_url = "https://www.myroms.org/svn/omlab/branches/arango" ;
		:svn_rev = "1124M" ;
		:code_dir = "/home/julia/ROMS/espresso/svn" ;
		:header_dir = "/home/julia/ROMS/espresso/Forward" ;
		:header_file = "espresso.h" ;
		:os = "Linux" ;
		:cpu = "x86_64" ;
		:compiler_system = "pgi" ;
		:compiler_command = "/opt/pgisoft/openmpi/bin/mpif90" ;
		:compiler_flags = " -O3 -tp k8-64 -Mfree" ;
		:tiling = "004x002" ;
		:history = "Thu Mar  8 11:45:22 2012: ncks -d ocean_time,879,881 http://tashtego.marine.rutgers.edu:8080/thredds/dodsC/roms/espresso/2009_da/avg roms.nc\n",
			"ROMS/TOMS, Version 3.2, Thursday - March 8, 2012 -  2:09:35 AM" ;
		:ana_file = "ROMS/Functionals/ana_btflux.h, /home/julia/ROMS/espresso/Forward/ana_nudgcoef.h" ;
		:CPP_options = "MyCPP, ADD_FSOBC, ADD_M2OBC, ANA_BSFLUX, ANA_BTFLUX, ASSUMED_SHAPE, AVERAGES, AVERAGES_AKS, AVERAGES_AKT, AVERAGES_FLUXES, BULK_FLUXES, CURVGRID, DJ_GRADPS, DOUBLE_PRECISION, EAST_FSCHAPMAN, EAST_M2FLATHER, EAST_M3NUDGING, EAST_M3RADIATION, EAST_TNUDGING, EAST_TRADIATION, EMINUSP, FORWARD_WRITE, !FULL_GRID, GLS_MIXING, KANTHA_CLAYSON, M3CLIMATOLOGY, M3CLM_NUDGING, MASKING, MIX_GEO_TS, MIX_S_UV, MPI, NONLINEAR, NONLIN_EOS, NORTHERN_WALL, N2S2_HORAVG, OBSERVATIONS, POWER_LAW, PROFILE, K_GSCHEME, RAMP_TIDES, !RST_SINGLE, SALINITY, SOLAR_SOURCE, SOLVE3D, SOUTH_FSCHAPMAN, SOUTH_M2FLATHER, SOUTH_M3NUDGING, SOUTH_M3RADIATION, SOUTH_TNUDGING, SOUTH_TRADIATION, SPLINES, SSH_TIDES, TCLIMATOLOGY, TCLM_NUDGING, TS_A4HADVECTION, TS_A4VADVECTION, TS_DIF2, TS_PSOURCE, UV_ADV, UV_COR, UV_U3HADVECTION, UV_C4VADVECTION, UV_QDRAG, UV_PSOURCE, UV_TIDES, UV_VIS2, VAR_RHO_2D, VERIFICATION, WEST_FSCHAPMAN, WEST_M2FLATHER, WEST_M3NUDGING, WEST_M3RADIATION, WEST_TNUDGING, WEST_TRADIATION" ;
		:NCO = "4.0.7" ;
}
